module vsdl

pub struct Version {
	major byte
	minor byte
	patch byte
}