module vsdl

pub enum RWWhence {
	start
	current
	end
}