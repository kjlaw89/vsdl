module gl

struct GLContext {
mut:
	ptr voidptr
}