module ttf

pub enum FontHinting {
	normal
	light
	mono
	@none
}

pub enum FontStyle {
	normal
	bold
	italic
	underline
	strikethrough
}