module ttf

pub struct Font {
mut:
	ptr voidptr
}
