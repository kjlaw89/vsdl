module mixer

// placeholder