module vsdl

pub struct RWops {
mut:
	ptr     voidptr
}