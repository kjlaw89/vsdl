module system

pub enum PowerState {
	unknown
	on_battery
	no_battery
	charging
	charged
}
